// Provides Cosine Lookup for I = 160

module CosineLookup (
	input wire clock,
	input wire [8:0] addr1,
	input wire [8:0] addr2,
	output logic [31:0] res1,
	output logic [31:0] res2
);

logic [31:0] lookup [0:319];

//does this work because of some packed/unpacked shenanigans??
always @(posedge clock) begin
	res1 <= lookup[{addr1}]<<7;
	res2 <= lookup[{addr2}]<<7;
end

// res = 1/I * cos(pi * addr / I)
// need to make sure addr is in [0, 2I)
assign lookup[0] = 32'h00cccccc; // 0 0.00625
assign lookup[1] = 32'h00ccc2b1; // 1 0.0062487952530129055
assign lookup[2] = 32'h00cca461; // 2 0.006245181476504518
assign lookup[3] = 32'h00cc71de; // 3 0.006239160063654475
assign lookup[4] = 32'h00cc2b2d; // 4 0.00623073333583205
assign lookup[5] = 32'h00cbd057; // 5 0.006219904541701231
assign lookup[6] = 32'h00cb6163; // 6 0.006206677855968289
assign lookup[7] = 32'h00cade5c; // 7 0.006191058377772358
assign lookup[8] = 32'h00ca4750; // 8 0.006173052128719611
assign lookup[9] = 32'h00c99c4d; // 9 0.006152666050561822
assign lookup[10] = 32'h00c8dd65; // 10 0.0061299080025201905
assign lookup[11] = 32'h00c80aa9; // 11 0.006104786758255453
assign lookup[12] = 32'h00c72430; // 12 0.0060773120024854785
assign lookup[13] = 32'h00c62a0f; // 13 0.006047494327251624
assign lookup[14] = 32'h00c51c5f; // 14 0.006015345227835296
assign lookup[15] = 32'h00c3fb3b; // 15 0.005980877098326305
assign lookup[16] = 32'h00c2c6c0; // 16 0.00594410322684471
assign lookup[17] = 32'h00c17f0c; // 17 0.005905037790417988
assign lookup[18] = 32'h00c0243e; // 18 0.005863695849515526
assign lookup[19] = 32'h00beb67b; // 19 0.005820093342242523
assign lookup[20] = 32'h00bd35e5; // 20 0.005774247078195542
assign lookup[21] = 32'h00bba2a2; // 21 0.0057261747319821
assign lookup[22] = 32'h00b9fcdb; // 22 0.005675894836406759
assign lookup[23] = 32'h00b844b9; // 23 0.005623426775326385
assign lookup[24] = 32'h00b67a67; // 24 0.005568790776177299
assign lookup[25] = 32'h00b49e12; // 25 0.005512007902177219
assign lookup[26] = 32'h00b2afeb; // 26 0.005453100044204982
assign lookup[27] = 32'h00b0b020; // 27 0.005392089912361199
assign lookup[28] = 32'h00ae9ee6; // 28 0.005329001027213077
assign lookup[29] = 32'h00ac7c70; // 29 0.005263857710726791
assign lookup[30] = 32'h00aa48f4; // 30 0.005196685076890908
assign lookup[31] = 32'h00a804a9; // 31 0.00512750902203446
assign lookup[32] = 32'h00a5afca; // 32 0.005056356214843421
assign lookup[33] = 32'h00a34a90; // 33 0.004983254086079419
assign lookup[34] = 32'h00a0d539; // 34 0.004908230818004656
assign lookup[35] = 32'h009e5002; // 35 0.004831315333517106
assign lookup[36] = 32'h009bbb2c; // 36 0.004752537285000193
assign lookup[37] = 32'h009916f6; // 37 0.00467192704289123
assign lookup[38] = 32'h009663a5; // 38 0.004589515683973035
assign lookup[39] = 32'h0093a17d; // 39 0.0045053349793932424
assign lookup[40] = 32'h0090d0c2; // 40 0.004419417382415922
assign lookup[41] = 32'h008df1bd; // 41 0.004331796015910225
assign lookup[42] = 32'h008b04b5; // 42 0.004242504659580886
assign lookup[43] = 32'h008809f5; // 43 0.004151577736945511
assign lookup[44] = 32'h008501c8; // 44 0.004059050302063648
assign lookup[45] = 32'h0081ec7a; // 45 0.003964958026022784
assign lookup[46] = 32'h007eca5a; // 46 0.003869337183186462
assign lookup[47] = 32'h007b9bb6; // 47 0.0037722246372098207
assign lookup[48] = 32'h007860e0; // 48 0.003673657826827957
assign lookup[49] = 32'h00751a28; // 49 0.003573674751422577
assign lookup[50] = 32'h0071c7e1; // 50 0.0034723139563725145
assign lookup[51] = 32'h006e6a60; // 51 0.0033696145181937526
assign lookup[52] = 32'h006b01f9; // 52 0.0032656160294746808
assign lookup[53] = 32'h00678f02; // 53 0.0031603585836124035
assign lookup[54] = 32'h006411d3; // 54 0.0030538827593559687
assign lookup[55] = 32'h00608ac3; // 55 0.002946229605162485
assign lookup[56] = 32'h005cfa2d; // 56 0.0028374406233721674
assign lookup[57] = 32'h00596069; // 57 0.0027275577542083887
assign lookup[58] = 32'h0055bdd3; // 58 0.0026166233596089257
assign lookup[59] = 32'h005212c7; // 59 0.0025046802068946316
assign lookup[60] = 32'h004e5fa2; // 60 0.0023917714522818114
assign lookup[61] = 32'h004aa4c0; // 61 0.002277940624244685
assign lookup[62] = 32'h0046e280; // 62 0.0021632316067343314
assign lookup[63] = 32'h00431941; // 63 0.002047688622260584
assign lookup[64] = 32'h003f4963; // 64 0.0019313562148434217
assign lookup[65] = 32'h003b7346; // 65 0.0018142792328403907
assign lookup[66] = 32'h0037974c; // 66 0.0016965028116567144
assign lookup[67] = 32'h0033b5d4; // 67 0.0015780723563447382
assign lookup[68] = 32'h002fcf42; // 68 0.0014590335240994093
assign lookup[69] = 32'h002be3f8; // 69 0.0013394322066565669
assign lookup[70] = 32'h0027f459; // 70 0.001219314512600802
assign lookup[71] = 32'h002400c9; // 71 0.0010987267495897153
assign lookup[72] = 32'h002009ab; // 72 0.0009777154065014433
assign lookup[73] = 32'h001c0f64; // 73 0.0008563271355123013
assign lookup[74] = 32'h00181258; // 74 0.0007346087341114857
assign lookup[75] = 32'h001412eb; // 75 0.0006126071270597548
assign lookup[76] = 32'h00101184; // 76 0.0004903693482990313
assign lookup[77] = 32'h000c0e86; // 77 0.00036794252281993113
assign lookup[78] = 32'h00080a58; // 78 0.00024537384849417917
assign lookup[79] = 32'h0004055e; // 79 0.00012271057787892656
assign lookup[80] = 32'h00000000; // 80 3.827021247335479e-19
assign lookup[81] = 32'hfffbfaa1; // 81 -0.0001227105778789258
assign lookup[82] = 32'hfff7f5a7; // 82 -0.00024537384849417706
assign lookup[83] = 32'hfff3f179; // 83 -0.0003679425228199318
assign lookup[84] = 32'hffefee7b; // 84 -0.0004903693482990305
assign lookup[85] = 32'hffebed14; // 85 -0.000612607127059754
assign lookup[86] = 32'hffe7eda7; // 86 -0.0007346087341114848
assign lookup[87] = 32'hffe3f09b; // 87 -0.0008563271355122991
assign lookup[88] = 32'hffdff654; // 88 -0.0009777154065014411
assign lookup[89] = 32'hffdbff36; // 89 -0.0010987267495897158
assign lookup[90] = 32'hffd80ba6; // 90 -0.0012193145126008012
assign lookup[91] = 32'hffd41c07; // 91 -0.0013394322066565662
assign lookup[92] = 32'hffd030bd; // 92 -0.0014590335240994084
assign lookup[93] = 32'hffcc4a2b; // 93 -0.001578072356344736
assign lookup[94] = 32'hffc868b3; // 94 -0.0016965028116567148
assign lookup[95] = 32'hffc48cb9; // 95 -0.00181427923284039
assign lookup[96] = 32'hffc0b69c; // 96 -0.0019313562148434208
assign lookup[97] = 32'hffbce6be; // 97 -0.002047688622260583
assign lookup[98] = 32'hffb91d7f; // 98 -0.0021632316067343293
assign lookup[99] = 32'hffb55b3f; // 99 -0.0022779406242446855
assign lookup[100] = 32'hffb1a05d; // 100 -0.002391771452281811
assign lookup[101] = 32'hffaded38; // 101 -0.002504680206894631
assign lookup[102] = 32'hffaa422c; // 102 -0.0026166233596089236
assign lookup[103] = 32'hffa69f96; // 103 -0.002727557754208387
assign lookup[104] = 32'hffa305d2; // 104 -0.0028374406233721674
assign lookup[105] = 32'hff9f753c; // 105 -0.0029462296051624855
assign lookup[106] = 32'hff9bee2c; // 106 -0.003053882759355969
assign lookup[107] = 32'hff9870fd; // 107 -0.0031603585836124026
assign lookup[108] = 32'hff94fe06; // 108 -0.00326561602947468
assign lookup[109] = 32'hff91959f; // 109 -0.003369614518193749
assign lookup[110] = 32'hff8e381e; // 110 -0.0034723139563725145
assign lookup[111] = 32'hff8ae5d7; // 111 -0.003573674751422576
assign lookup[112] = 32'hff879f1f; // 112 -0.0036736578268279562
assign lookup[113] = 32'hff846449; // 113 -0.0037722246372098216
assign lookup[114] = 32'hff8135a5; // 114 -0.003869337183186461
assign lookup[115] = 32'hff7e1385; // 115 -0.003964958026022786
assign lookup[116] = 32'hff7afe37; // 116 -0.004059050302063647
assign lookup[117] = 32'hff77f60a; // 117 -0.004151577736945511
assign lookup[118] = 32'hff74fb4a; // 118 -0.004242504659580884
assign lookup[119] = 32'hff720e42; // 119 -0.004331796015910223
assign lookup[120] = 32'hff6f2f3d; // 120 -0.004419417382415922
assign lookup[121] = 32'hff6c5e82; // 121 -0.0045053349793932424
assign lookup[122] = 32'hff699c5a; // 122 -0.004589515683973035
assign lookup[123] = 32'hff66e909; // 123 -0.004671927042891229
assign lookup[124] = 32'hff6444d3; // 124 -0.004752537285000193
assign lookup[125] = 32'hff61affd; // 125 -0.004831315333517104
assign lookup[126] = 32'hff5f2ac6; // 126 -0.004908230818004656
assign lookup[127] = 32'hff5cb56f; // 127 -0.004983254086079419
assign lookup[128] = 32'hff5a5035; // 128 -0.0050563562148434205
assign lookup[129] = 32'hff57fb56; // 129 -0.00512750902203446
assign lookup[130] = 32'hff55b70b; // 130 -0.005196685076890906
assign lookup[131] = 32'hff53838f; // 131 -0.005263857710726792
assign lookup[132] = 32'hff516119; // 132 -0.005329001027213076
assign lookup[133] = 32'hff4f4fdf; // 133 -0.005392089912361199
assign lookup[134] = 32'hff4d5014; // 134 -0.005453100044204981
assign lookup[135] = 32'hff4b61ed; // 135 -0.0055120079021772185
assign lookup[136] = 32'hff498598; // 136 -0.005568790776177298
assign lookup[137] = 32'hff47bb46; // 137 -0.005623426775326384
assign lookup[138] = 32'hff460324; // 138 -0.005675894836406759
assign lookup[139] = 32'hff445d5d; // 139 -0.005726174731982099
assign lookup[140] = 32'hff42ca1a; // 140 -0.005774247078195542
assign lookup[141] = 32'hff414984; // 141 -0.005820093342242521
assign lookup[142] = 32'hff3fdbc1; // 142 -0.005863695849515526
assign lookup[143] = 32'hff3e80f3; // 143 -0.005905037790417987
assign lookup[144] = 32'hff3d393f; // 144 -0.00594410322684471
assign lookup[145] = 32'hff3c04c4; // 145 -0.005980877098326305
assign lookup[146] = 32'hff3ae3a0; // 146 -0.006015345227835295
assign lookup[147] = 32'hff39d5f0; // 147 -0.006047494327251624
assign lookup[148] = 32'hff38dbcf; // 148 -0.0060773120024854785
assign lookup[149] = 32'hff37f556; // 149 -0.006104786758255452
assign lookup[150] = 32'hff37229a; // 150 -0.0061299080025201905
assign lookup[151] = 32'hff3663b2; // 151 -0.006152666050561822
assign lookup[152] = 32'hff35b8af; // 152 -0.0061730521287196105
assign lookup[153] = 32'hff3521a3; // 153 -0.006191058377772358
assign lookup[154] = 32'hff349e9c; // 154 -0.006206677855968289
assign lookup[155] = 32'hff342fa8; // 155 -0.00621990454170123
assign lookup[156] = 32'hff33d4d2; // 156 -0.00623073333583205
assign lookup[157] = 32'hff338e21; // 157 -0.006239160063654474
assign lookup[158] = 32'hff335b9e; // 158 -0.006245181476504518
assign lookup[159] = 32'hff333d4e; // 159 -0.0062487952530129055
assign lookup[160] = 32'hff333333; // 160 -0.00625
assign lookup[161] = 32'hff333d4e; // 161 -0.0062487952530129055
assign lookup[162] = 32'hff335b9e; // 162 -0.006245181476504518
assign lookup[163] = 32'hff338e21; // 163 -0.006239160063654475
assign lookup[164] = 32'hff33d4d2; // 164 -0.00623073333583205
assign lookup[165] = 32'hff342fa8; // 165 -0.006219904541701231
assign lookup[166] = 32'hff349e9c; // 166 -0.006206677855968289
assign lookup[167] = 32'hff3521a3; // 167 -0.006191058377772358
assign lookup[168] = 32'hff35b8af; // 168 -0.006173052128719611
assign lookup[169] = 32'hff3663b2; // 169 -0.006152666050561822
assign lookup[170] = 32'hff37229a; // 170 -0.0061299080025201905
assign lookup[171] = 32'hff37f556; // 171 -0.006104786758255453
assign lookup[172] = 32'hff38dbcf; // 172 -0.006077312002485479
assign lookup[173] = 32'hff39d5f0; // 173 -0.006047494327251624
assign lookup[174] = 32'hff3ae3a0; // 174 -0.006015345227835296
assign lookup[175] = 32'hff3c04c4; // 175 -0.005980877098326306
assign lookup[176] = 32'hff3d393f; // 176 -0.005944103226844711
assign lookup[177] = 32'hff3e80f3; // 177 -0.005905037790417988
assign lookup[178] = 32'hff3fdbc1; // 178 -0.005863695849515526
assign lookup[179] = 32'hff414984; // 179 -0.005820093342242522
assign lookup[180] = 32'hff42ca1a; // 180 -0.005774247078195543
assign lookup[181] = 32'hff445d5d; // 181 -0.0057261747319821
assign lookup[182] = 32'hff460324; // 182 -0.005675894836406759
assign lookup[183] = 32'hff47bb46; // 183 -0.0056234267753263855
assign lookup[184] = 32'hff498598; // 184 -0.005568790776177299
assign lookup[185] = 32'hff4b61ed; // 185 -0.00551200790217722
assign lookup[186] = 32'hff4d5014; // 186 -0.005453100044204983
assign lookup[187] = 32'hff4f4fdf; // 187 -0.005392089912361198
assign lookup[188] = 32'hff516119; // 188 -0.005329001027213075
assign lookup[189] = 32'hff53838f; // 189 -0.005263857710726791
assign lookup[190] = 32'hff55b70b; // 190 -0.005196685076890908
assign lookup[191] = 32'hff57fb56; // 191 -0.005127509022034462
assign lookup[192] = 32'hff5a5035; // 192 -0.005056356214843421
assign lookup[193] = 32'hff5cb56f; // 193 -0.004983254086079419
assign lookup[194] = 32'hff5f2ac6; // 194 -0.0049082308180046575
assign lookup[195] = 32'hff61affd; // 195 -0.004831315333517107
assign lookup[196] = 32'hff6444d3; // 196 -0.0047525372850001964
assign lookup[197] = 32'hff66e909; // 197 -0.0046719270428912316
assign lookup[198] = 32'hff699c5a; // 198 -0.004589515683973035
assign lookup[199] = 32'hff6c5e82; // 199 -0.004505334979393242
assign lookup[200] = 32'hff6f2f3d; // 200 -0.004419417382415923
assign lookup[201] = 32'hff720e42; // 201 -0.004331796015910224
assign lookup[202] = 32'hff74fb4a; // 202 -0.004242504659580886
assign lookup[203] = 32'hff77f60a; // 203 -0.0041515777369455125
assign lookup[204] = 32'hff7afe37; // 204 -0.004059050302063651
assign lookup[205] = 32'hff7e1385; // 205 -0.003964958026022787
assign lookup[206] = 32'hff8135a5; // 206 -0.0038693371831864643
assign lookup[207] = 32'hff846449; // 207 -0.003772224637209823
assign lookup[208] = 32'hff879f1f; // 208 -0.003673657826827958
assign lookup[209] = 32'hff8ae5d7; // 209 -0.003573674751422577
assign lookup[210] = 32'hff8e381e; // 210 -0.0034723139563725136
assign lookup[211] = 32'hff91959f; // 211 -0.0033696145181937504
assign lookup[212] = 32'hff94fe06; // 212 -0.0032656160294746786
assign lookup[213] = 32'hff9870fd; // 213 -0.003160358583612406
assign lookup[214] = 32'hff9bee2c; // 214 -0.0030538827593559704
assign lookup[215] = 32'hff9f753c; // 215 -0.002946229605162487
assign lookup[216] = 32'hffa305d2; // 216 -0.0028374406233721682
assign lookup[217] = 32'hffa69f96; // 217 -0.0027275577542083883
assign lookup[218] = 32'hffaa422c; // 218 -0.0026166233596089305
assign lookup[219] = 32'hffaded38; // 219 -0.00250468020689463
assign lookup[220] = 32'hffb1a05d; // 220 -0.0023917714522818092
assign lookup[221] = 32'hffb55b3f; // 221 -0.0022779406242446833
assign lookup[222] = 32'hffb91d7f; // 222 -0.0021632316067343336
assign lookup[223] = 32'hffbce6be; // 223 -0.002047688622260586
assign lookup[224] = 32'hffc0b69c; // 224 -0.0019313562148434223
assign lookup[225] = 32'hffc48cb9; // 225 -0.0018142792328403902
assign lookup[226] = 32'hffc868b3; // 226 -0.0016965028116567138
assign lookup[227] = 32'hffcc4a2b; // 227 -0.0015780723563447417
assign lookup[228] = 32'hffd030bd; // 228 -0.0014590335240994125
assign lookup[229] = 32'hffd41c07; // 229 -0.0013394322066565703
assign lookup[230] = 32'hffd80ba6; // 230 -0.0012193145126007986
assign lookup[231] = 32'hffdbff36; // 231 -0.0010987267495897175
assign lookup[232] = 32'hffdff654; // 232 -0.000977715406501444
assign lookup[233] = 32'hffe3f09b; // 233 -0.0008563271355123006
assign lookup[234] = 32'hffe7eda7; // 234 -0.000734608734111485
assign lookup[235] = 32'hffebed14; // 235 -0.0006126071270597528
assign lookup[236] = 32'hffefee7b; // 236 -0.0004903693482990348
assign lookup[237] = 32'hfff3f179; // 237 -0.00036794252281993465
assign lookup[238] = 32'hfff7f5a7; // 238 -0.00024537384849418134
assign lookup[239] = 32'hfffbfaa1; // 239 -0.00012271057787892873
assign lookup[240] = 32'h00000000; // 240 -1.1481063742006436e-18
assign lookup[241] = 32'h0004055e; // 241 0.00012271057787892643
assign lookup[242] = 32'h00080a58; // 242 0.000245373848494179
assign lookup[243] = 32'h000c0e86; // 243 0.0003679425228199324
assign lookup[244] = 32'h00101184; // 244 0.0004903693482990326
assign lookup[245] = 32'h001412eb; // 245 0.0006126071270597506
assign lookup[246] = 32'h00181258; // 246 0.0007346087341114827
assign lookup[247] = 32'h001c0f64; // 247 0.0008563271355122984
assign lookup[248] = 32'h002009ab; // 248 0.0009777154065014418
assign lookup[249] = 32'h002400c9; // 249 0.0010987267495897151
assign lookup[250] = 32'h0027f459; // 250 0.0012193145126007964
assign lookup[251] = 32'h002be3f8; // 251 0.001339432206656568
assign lookup[252] = 32'h002fcf42; // 252 0.0014590335240994103
assign lookup[253] = 32'h0033b5d4; // 253 0.0015780723563447393
assign lookup[254] = 32'h0037974c; // 254 0.0016965028116567118
assign lookup[255] = 32'h003b7346; // 255 0.0018142792328403878
assign lookup[256] = 32'h003f4963; // 256 0.0019313562148434201
assign lookup[257] = 32'h00431941; // 257 0.002047688622260584
assign lookup[258] = 32'h0046e280; // 258 0.0021632316067343314
assign lookup[259] = 32'h004aa4c0; // 259 0.002277940624244681
assign lookup[260] = 32'h004e5fa2; // 260 0.0023917714522818075
assign lookup[261] = 32'h005212c7; // 261 0.0025046802068946277
assign lookup[262] = 32'h0055bdd3; // 262 0.0026166233596089284
assign lookup[263] = 32'h00596069; // 263 0.002727557754208386
assign lookup[264] = 32'h005cfa2d; // 264 0.0028374406233721665
assign lookup[265] = 32'h00608ac3; // 265 0.002946229605162485
assign lookup[266] = 32'h006411d3; // 266 0.0030538827593559687
assign lookup[267] = 32'h00678f02; // 267 0.0031603585836124043
assign lookup[268] = 32'h006b01f9; // 268 0.0032656160294746773
assign lookup[269] = 32'h006e6a60; // 269 0.0033696145181937483
assign lookup[270] = 32'h0071c7e1; // 270 0.0034723139563725114
assign lookup[271] = 32'h00751a28; // 271 0.003573674751422575
assign lookup[272] = 32'h007860e0; // 272 0.003673657826827956
assign lookup[273] = 32'h007b9bb6; // 273 0.0037722246372098207
assign lookup[274] = 32'h007eca5a; // 274 0.003869337183186462
assign lookup[275] = 32'h0081ec7a; // 275 0.003964958026022785
assign lookup[276] = 32'h008501c8; // 276 0.004059050302063649
assign lookup[277] = 32'h008809f5; // 277 0.004151577736945508
assign lookup[278] = 32'h008b04b5; // 278 0.004242504659580884
assign lookup[279] = 32'h008df1bd; // 279 0.0043317960159102225
assign lookup[280] = 32'h0090d0c2; // 280 0.004419417382415921
assign lookup[281] = 32'h0093a17d; // 281 0.004505334979393242
assign lookup[282] = 32'h009663a5; // 282 0.004589515683973031
assign lookup[283] = 32'h009916f6; // 283 0.00467192704289123
assign lookup[284] = 32'h009bbb2c; // 284 0.004752537285000194
assign lookup[285] = 32'h009e5002; // 285 0.004831315333517107
assign lookup[286] = 32'h00a0d539; // 286 0.004908230818004654
assign lookup[287] = 32'h00a34a90; // 287 0.004983254086079418
assign lookup[288] = 32'h00a5afca; // 288 0.0050563562148434205
assign lookup[289] = 32'h00a804a9; // 289 0.00512750902203446
assign lookup[290] = 32'h00aa48f4; // 290 0.005196685076890908
assign lookup[291] = 32'h00ac7c70; // 291 0.0052638577107267884
assign lookup[292] = 32'h00ae9ee6; // 292 0.005329001027213074
assign lookup[293] = 32'h00b0b020; // 293 0.005392089912361197
assign lookup[294] = 32'h00b2afeb; // 294 0.005453100044204983
assign lookup[295] = 32'h00b49e12; // 295 0.005512007902177218
assign lookup[296] = 32'h00b67a67; // 296 0.005568790776177298
assign lookup[297] = 32'h00b844b9; // 297 0.005623426775326384
assign lookup[298] = 32'h00b9fcdb; // 298 0.005675894836406758
assign lookup[299] = 32'h00bba2a2; // 299 0.0057261747319821
assign lookup[300] = 32'h00bd35e5; // 300 0.005774247078195541
assign lookup[301] = 32'h00beb67b; // 301 0.005820093342242521
assign lookup[302] = 32'h00c0243e; // 302 0.005863695849515524
assign lookup[303] = 32'h00c17f0c; // 303 0.005905037790417987
assign lookup[304] = 32'h00c2c6c0; // 304 0.00594410322684471
assign lookup[305] = 32'h00c3fb3b; // 305 0.005980877098326305
assign lookup[306] = 32'h00c51c5f; // 306 0.006015345227835296
assign lookup[307] = 32'h00c62a0f; // 307 0.006047494327251624
assign lookup[308] = 32'h00c72430; // 308 0.006077312002485479
assign lookup[309] = 32'h00c80aa9; // 309 0.0061047867582554515
assign lookup[310] = 32'h00c8dd65; // 310 0.00612990800252019
assign lookup[311] = 32'h00c99c4d; // 311 0.006152666050561822
assign lookup[312] = 32'h00ca4750; // 312 0.0061730521287196105
assign lookup[313] = 32'h00cade5c; // 313 0.006191058377772358
assign lookup[314] = 32'h00cb6163; // 314 0.006206677855968288
assign lookup[315] = 32'h00cbd057; // 315 0.006219904541701231
assign lookup[316] = 32'h00cc2b2d; // 316 0.00623073333583205
assign lookup[317] = 32'h00cc71de; // 317 0.006239160063654475
assign lookup[318] = 32'h00cca461; // 318 0.006245181476504518
assign lookup[319] = 32'h00ccc2b1; // 319 0.0062487952530129055

endmodule