// Provides hamming window factor for windowing step before fft.
// assumes 400 samples per window.

module Hamming (
	input clock,
	input [8:0] addr,
	output [31:0] hamming_factor
);

logic [31:0] ham [0:399];
logic [31:0] ham_register;

//does this work because of some packed/unpacked shenanigans??
always @(posedge clock) begin
	ham_register <= ham[{addr}];
end

assign hamming_factor = ham_register;

// table of hamming window values (just 1 for now.)
//      wn_re = 0.54 - 0.46*cos(-2pi*n/400)  
assign  ham[ 0] = 32'h00000000;   //  0  0.080 
assign  ham[ 1] = 32'h0A3F4CB0;   //  1  0.080 
assign  ham[ 2] = 32'h0A44E0B4;   //  2  0.080 
assign  ham[ 3] = 32'h0A4E2C59;   //  3  0.081 
assign  ham[ 4] = 32'h0A5B2F05;   //  4  0.081 
assign  ham[ 5] = 32'h0A6BE7E9;   //  5  0.081 
assign  ham[ 6] = 32'h0A8055F4;   //  6  0.082 
assign  ham[ 7] = 32'h0A9877DD;   //  7  0.083 
assign  ham[ 8] = 32'h0AB44C1D;   //  8  0.084 
assign  ham[ 9] = 32'h0AD3D0F3;   //  9  0.085 
assign  ham[10] = 32'h0AF70460;   // 10  0.086 
assign  ham[11] = 32'h0B1DE42C;   // 11  0.087 
assign  ham[12] = 32'h0B486DE2;   // 12  0.088 
assign  ham[13] = 32'h0B769ED2;   // 13  0.090 
assign  ham[14] = 32'h0BA87411;   // 14  0.091 
assign  ham[15] = 32'h0BDDEA7A;   // 15  0.093 
assign  ham[16] = 32'h0C16FEAC;   // 16  0.094 
assign  ham[17] = 32'h0C53AD0B;   // 17  0.096 
assign  ham[18] = 32'h0C93F1C4;   // 18  0.098 
assign  ham[19] = 32'h0CD7C8C6;   // 19  0.100 
assign  ham[20] = 32'h0D1F2DC8;   // 20  0.103 
assign  ham[21] = 32'h0D6A1C49;   // 21  0.105 
assign  ham[22] = 32'h0DB88F8C;   // 22  0.107 
assign  ham[23] = 32'h0E0A829C;   // 23  0.110 
assign  ham[24] = 32'h0E5FF04E;   // 24  0.112 
assign  ham[25] = 32'h0EB8D33B;   // 25  0.115 
assign  ham[26] = 32'h0F1525C6;   // 26  0.118 
assign  ham[27] = 32'h0F74E21B;   // 27  0.121 
assign  ham[28] = 32'h0FD8022C;   // 28  0.124 
assign  ham[29] = 32'h103E7FB8;   // 29  0.127 
assign  ham[30] = 32'h10A85445;   // 30  0.130 
assign  ham[31] = 32'h11157924;   // 31  0.133 
assign  ham[32] = 32'h1185E770;   // 32  0.137 
assign  ham[33] = 32'h11F9980E;   // 33  0.140 
assign  ham[34] = 32'h127083B1;   // 34  0.144 
assign  ham[35] = 32'h12EAA2D5;   // 35  0.148 
assign  ham[36] = 32'h1367EDC4;   // 36  0.152 
assign  ham[37] = 32'h13E85C93;   // 37  0.156 
assign  ham[38] = 32'h146BE726;   // 38  0.160 
assign  ham[39] = 32'h14F2852E;   // 39  0.164 
assign  ham[40] = 32'h157C2E29;   // 40  0.168 
assign  ham[41] = 32'h1608D967;   // 41  0.172 
assign  ham[42] = 32'h16987E04;   // 42  0.177 
assign  ham[43] = 32'h172B12EE;   // 43  0.181 
assign  ham[44] = 32'h17C08EE3;   // 44  0.186 
assign  ham[45] = 32'h1858E871;   // 45  0.190 
assign  ham[46] = 32'h18F415F8;   // 46  0.195 
assign  ham[47] = 32'h19920DAC;   // 47  0.200 
assign  ham[48] = 32'h1A32C593;   // 48  0.205 
assign  ham[49] = 32'h1AD63384;   // 49  0.210 
assign  ham[50] = 32'h1B7C4D2F;   // 50  0.215 
assign  ham[51] = 32'h1C250814;   // 51  0.220 
assign  ham[52] = 32'h1CD0598C;   // 52  0.225 
assign  ham[53] = 32'h1D7E36C5;   // 53  0.230 
assign  ham[54] = 32'h1E2E94C2;   // 54  0.236 
assign  ham[55] = 32'h1EE16860;   // 55  0.241 
assign  ham[56] = 32'h1F96A654;   // 56  0.247 
assign  ham[57] = 32'h204E432B;   // 57  0.252 
assign  ham[58] = 32'h2108334B;   // 58  0.258 
assign  ham[59] = 32'h21C46AF7;   // 59  0.264 
assign  ham[60] = 32'h2282DE4A;   // 60  0.270 
assign  ham[61] = 32'h2343813D;   // 61  0.275 
assign  ham[62] = 32'h240647A5;   // 62  0.281 
assign  ham[63] = 32'h24CB2535;   // 63  0.287 
assign  ham[64] = 32'h25920D7D;   // 64  0.294 
assign  ham[65] = 32'h265AF3ED;   // 65  0.300 
assign  ham[66] = 32'h2725CBD4;   // 66  0.306 
assign  ham[67] = 32'h27F28863;   // 67  0.312 
assign  ham[68] = 32'h28C11CAB;   // 68  0.318 
assign  ham[69] = 32'h29917B9F;   // 69  0.325 
assign  ham[70] = 32'h2A639816;   // 70  0.331 
assign  ham[71] = 32'h2B3764CA;   // 71  0.338 
assign  ham[72] = 32'h2C0CD45B;   // 72  0.344 
assign  ham[73] = 32'h2CE3D94E;   // 73  0.351 
assign  ham[74] = 32'h2DBC660D;   // 74  0.357 
assign  ham[75] = 32'h2E966CEC;   // 75  0.364 
assign  ham[76] = 32'h2F71E024;   // 76  0.371 
assign  ham[77] = 32'h304EB1D8;   // 77  0.377 
assign  ham[78] = 32'h312CD417;   // 78  0.384 
assign  ham[79] = 32'h320C38D9;   // 79  0.391 
assign  ham[80] = 32'h32ECD200;   // 80  0.398 
assign  ham[81] = 32'h33CE915E;   // 81  0.405 
assign  ham[82] = 32'h34B168B0;   // 82  0.412 
assign  ham[83] = 32'h359549A2;   // 83  0.419 
assign  ham[84] = 32'h367A25D0;   // 84  0.426 
assign  ham[85] = 32'h375FEEC3;   // 85  0.433 
assign  ham[86] = 32'h384695FA;   // 86  0.440 
assign  ham[87] = 32'h392E0CE2;   // 87  0.447 
assign  ham[88] = 32'h3A1644DC;   // 88  0.454 
assign  ham[89] = 32'h3AFF2F3D;   // 89  0.461 
assign  ham[90] = 32'h3BE8BD50;   // 90  0.468 
assign  ham[91] = 32'h3CD2E054;   // 91  0.475 
assign  ham[92] = 32'h3DBD897E;   // 92  0.482 
assign  ham[93] = 32'h3EA8A9FC;   // 93  0.490 
assign  ham[94] = 32'h3F9432F4;   // 94  0.497 
assign  ham[95] = 32'h40801586;   // 95  0.504 
assign  ham[96] = 32'h416C42CC;   // 96  0.511 
assign  ham[97] = 32'h4258ABD9;   // 97  0.518 
assign  ham[98] = 32'h434541C0;   // 98  0.526 
assign  ham[99] = 32'h4431F58F;   // 99  0.533 
assign  ham[100] = 32'h451EB852;   // 100  0.540 
assign  ham[101] = 32'h460B7B15;   // 101  0.547 
assign  ham[102] = 32'h46F82EE4;   // 102  0.554 
assign  ham[103] = 32'h47E4C4CB;   // 103  0.562 
assign  ham[104] = 32'h48D12DD8;   // 104  0.569 
assign  ham[105] = 32'h49BD5B1D;   // 105  0.576 
assign  ham[106] = 32'h4AA93DAF;   // 106  0.583 
assign  ham[107] = 32'h4B94C6A8;   // 107  0.590 
assign  ham[108] = 32'h4C7FE726;   // 108  0.598 
assign  ham[109] = 32'h4D6A9050;   // 109  0.605 
assign  ham[110] = 32'h4E54B354;   // 110  0.612 
assign  ham[111] = 32'h4F3E4166;   // 111  0.619 
assign  ham[112] = 32'h50272BC8;   // 112  0.626 
assign  ham[113] = 32'h510F63C2;   // 113  0.633 
assign  ham[114] = 32'h51F6DAAA;   // 114  0.640 
assign  ham[115] = 32'h52DD81E1;   // 115  0.647 
assign  ham[116] = 32'h53C34AD4;   // 116  0.654 
assign  ham[117] = 32'h54A82701;   // 117  0.661 
assign  ham[118] = 32'h558C07F3;   // 118  0.668 
assign  ham[119] = 32'h566EDF45;   // 119  0.675 
assign  ham[120] = 32'h57509EA3;   // 120  0.682 
assign  ham[121] = 32'h583137CB;   // 121  0.689 
assign  ham[122] = 32'h59109C8C;   // 122  0.696 
assign  ham[123] = 32'h59EEBECC;   // 123  0.703 
assign  ham[124] = 32'h5ACB9080;   // 124  0.709 
assign  ham[125] = 32'h5BA703B8;   // 125  0.716 
assign  ham[126] = 32'h5C810A96;   // 126  0.723 
assign  ham[127] = 32'h5D599756;   // 127  0.729 
assign  ham[128] = 32'h5E309C48;   // 128  0.736 
assign  ham[129] = 32'h5F060BDA;   // 129  0.742 
assign  ham[130] = 32'h5FD9D88E;   // 130  0.749 
assign  ham[131] = 32'h60ABF505;   // 131  0.755 
assign  ham[132] = 32'h617C53F9;   // 132  0.762 
assign  ham[133] = 32'h624AE841;   // 133  0.768 
assign  ham[134] = 32'h6317A4D0;   // 134  0.774 
assign  ham[135] = 32'h63E27CB7;   // 135  0.780 
assign  ham[136] = 32'h64AB6327;   // 136  0.786 
assign  ham[137] = 32'h65724B6F;   // 137  0.793 
assign  ham[138] = 32'h663728FF;   // 138  0.799 
assign  ham[139] = 32'h66F9EF67;   // 139  0.805 
assign  ham[140] = 32'h67BA925A;   // 140  0.810 
assign  ham[141] = 32'h687905AD;   // 141  0.816 
assign  ham[142] = 32'h69353D59;   // 142  0.822 
assign  ham[143] = 32'h69EF2D79;   // 143  0.828 
assign  ham[144] = 32'h6AA6CA50;   // 144  0.833 
assign  ham[145] = 32'h6B5C0843;   // 145  0.839 
assign  ham[146] = 32'h6C0EDBE2;   // 146  0.844 
assign  ham[147] = 32'h6CBF39DF;   // 147  0.850 
assign  ham[148] = 32'h6D6D1717;   // 148  0.855 
assign  ham[149] = 32'h6E18688F;   // 149  0.860 
assign  ham[150] = 32'h6EC12375;   // 150  0.865 
assign  ham[151] = 32'h6F673D1F;   // 151  0.870 
assign  ham[152] = 32'h700AAB11;   // 152  0.875 
assign  ham[153] = 32'h70AB62F8;   // 153  0.880 
assign  ham[154] = 32'h71495AAC;   // 154  0.885 
assign  ham[155] = 32'h71E48833;   // 155  0.890 
assign  ham[156] = 32'h727CE1C1;   // 156  0.894 
assign  ham[157] = 32'h73125DB5;   // 157  0.899 
assign  ham[158] = 32'h73A4F29F;   // 158  0.903 
assign  ham[159] = 32'h7434973D;   // 159  0.908 
assign  ham[160] = 32'h74C1427A;   // 160  0.912 
assign  ham[161] = 32'h754AEB76;   // 161  0.916 
assign  ham[162] = 32'h75D1897E;   // 162  0.920 
assign  ham[163] = 32'h76551411;   // 163  0.924 
assign  ham[164] = 32'h76D582E0;   // 164  0.928 
assign  ham[165] = 32'h7752CDCF;   // 165  0.932 
assign  ham[166] = 32'h77CCECF3;   // 166  0.936 
assign  ham[167] = 32'h7843D896;   // 167  0.940 
assign  ham[168] = 32'h78B78934;   // 168  0.943 
assign  ham[169] = 32'h7927F780;   // 169  0.947 
assign  ham[170] = 32'h79951C5F;   // 170  0.950 
assign  ham[171] = 32'h79FEF0EC;   // 171  0.953 
assign  ham[172] = 32'h7A656E78;   // 172  0.956 
assign  ham[173] = 32'h7AC88E89;   // 173  0.959 
assign  ham[174] = 32'h7B284ADE;   // 174  0.962 
assign  ham[175] = 32'h7B849D69;   // 175  0.965 
assign  ham[176] = 32'h7BDD8056;   // 176  0.968 
assign  ham[177] = 32'h7C32EE07;   // 177  0.970 
assign  ham[178] = 32'h7C84E118;   // 178  0.973 
assign  ham[179] = 32'h7CD3545B;   // 179  0.975 
assign  ham[180] = 32'h7D1E42DC;   // 180  0.977 
assign  ham[181] = 32'h7D65A7DE;   // 181  0.980 
assign  ham[182] = 32'h7DA97EE0;   // 182  0.982 
assign  ham[183] = 32'h7DE9C398;   // 183  0.984 
assign  ham[184] = 32'h7E2671F8;   // 184  0.986 
assign  ham[185] = 32'h7E5F862A;   // 185  0.987 
assign  ham[186] = 32'h7E94FC92;   // 186  0.989 
assign  ham[187] = 32'h7EC6D1D2;   // 187  0.990 
assign  ham[188] = 32'h7EF502C2;   // 188  0.992 
assign  ham[189] = 32'h7F1F8C78;   // 189  0.993 
assign  ham[190] = 32'h7F466C44;   // 190  0.994 
assign  ham[191] = 32'h7F699FB1;   // 191  0.995 
assign  ham[192] = 32'h7F892487;   // 192  0.996 
assign  ham[193] = 32'h7FA4F8C7;   // 193  0.997 
assign  ham[194] = 32'h7FBD1AB0;   // 194  0.998 
assign  ham[195] = 32'h7FD188BB;   // 195  0.999 
assign  ham[196] = 32'h7FE2419F;   // 196  0.999 
assign  ham[197] = 32'h7FEF444B;   // 197  0.999 
assign  ham[198] = 32'h7FF88FEF;   // 198  1.000 
assign  ham[199] = 32'h7FFE23F4;   // 199  1.000 
assign  ham[200] = 32'h7FFFFFFF;   // 200  1.000 
assign  ham[201] = 32'h7FFE23F4;   // 201  1.000 
assign  ham[202] = 32'h7FF88FEF;   // 202  1.000 
assign  ham[203] = 32'h7FEF444B;   // 203  0.999 
assign  ham[204] = 32'h7FE2419F;   // 204  0.999 
assign  ham[205] = 32'h7FD188BB;   // 205  0.999 
assign  ham[206] = 32'h7FBD1AB0;   // 206  0.998 
assign  ham[207] = 32'h7FA4F8C7;   // 207  0.997 
assign  ham[208] = 32'h7F892487;   // 208  0.996 
assign  ham[209] = 32'h7F699FB1;   // 209  0.995 
assign  ham[210] = 32'h7F466C44;   // 210  0.994 
assign  ham[211] = 32'h7F1F8C78;   // 211  0.993 
assign  ham[212] = 32'h7EF502C2;   // 212  0.992 
assign  ham[213] = 32'h7EC6D1D2;   // 213  0.990 
assign  ham[214] = 32'h7E94FC92;   // 214  0.989 
assign  ham[215] = 32'h7E5F862A;   // 215  0.987 
assign  ham[216] = 32'h7E2671F8;   // 216  0.986 
assign  ham[217] = 32'h7DE9C398;   // 217  0.984 
assign  ham[218] = 32'h7DA97EE0;   // 218  0.982 
assign  ham[219] = 32'h7D65A7DE;   // 219  0.980 
assign  ham[220] = 32'h7D1E42DC;   // 220  0.977 
assign  ham[221] = 32'h7CD3545B;   // 221  0.975 
assign  ham[222] = 32'h7C84E118;   // 222  0.973 
assign  ham[223] = 32'h7C32EE07;   // 223  0.970 
assign  ham[224] = 32'h7BDD8056;   // 224  0.968 
assign  ham[225] = 32'h7B849D69;   // 225  0.965 
assign  ham[226] = 32'h7B284ADE;   // 226  0.962 
assign  ham[227] = 32'h7AC88E89;   // 227  0.959 
assign  ham[228] = 32'h7A656E78;   // 228  0.956 
assign  ham[229] = 32'h79FEF0EC;   // 229  0.953 
assign  ham[230] = 32'h79951C5F;   // 230  0.950 
assign  ham[231] = 32'h7927F780;   // 231  0.947 
assign  ham[232] = 32'h78B78934;   // 232  0.943 
assign  ham[233] = 32'h7843D896;   // 233  0.940 
assign  ham[234] = 32'h77CCECF3;   // 234  0.936 
assign  ham[235] = 32'h7752CDCF;   // 235  0.932 
assign  ham[236] = 32'h76D582E0;   // 236  0.928 
assign  ham[237] = 32'h76551411;   // 237  0.924 
assign  ham[238] = 32'h75D1897E;   // 238  0.920 
assign  ham[239] = 32'h754AEB76;   // 239  0.916 
assign  ham[240] = 32'h74C1427A;   // 240  0.912 
assign  ham[241] = 32'h7434973D;   // 241  0.908 
assign  ham[242] = 32'h73A4F29F;   // 242  0.903 
assign  ham[243] = 32'h73125DB5;   // 243  0.899 
assign  ham[244] = 32'h727CE1C1;   // 244  0.894 
assign  ham[245] = 32'h71E48833;   // 245  0.890 
assign  ham[246] = 32'h71495AAC;   // 246  0.885 
assign  ham[247] = 32'h70AB62F8;   // 247  0.880 
assign  ham[248] = 32'h700AAB11;   // 248  0.875 
assign  ham[249] = 32'h6F673D1F;   // 249  0.870 
assign  ham[250] = 32'h6EC12375;   // 250  0.865 
assign  ham[251] = 32'h6E18688F;   // 251  0.860 
assign  ham[252] = 32'h6D6D1717;   // 252  0.855 
assign  ham[253] = 32'h6CBF39DF;   // 253  0.850 
assign  ham[254] = 32'h6C0EDBE2;   // 254  0.844 
assign  ham[255] = 32'h6B5C0843;   // 255  0.839 
assign  ham[256] = 32'h6AA6CA50;   // 256  0.833 
assign  ham[257] = 32'h69EF2D79;   // 257  0.828 
assign  ham[258] = 32'h69353D59;   // 258  0.822 
assign  ham[259] = 32'h687905AD;   // 259  0.816 
assign  ham[260] = 32'h67BA925A;   // 260  0.810 
assign  ham[261] = 32'h66F9EF67;   // 261  0.805 
assign  ham[262] = 32'h663728FF;   // 262  0.799 
assign  ham[263] = 32'h65724B6F;   // 263  0.793 
assign  ham[264] = 32'h64AB6327;   // 264  0.786 
assign  ham[265] = 32'h63E27CB7;   // 265  0.780 
assign  ham[266] = 32'h6317A4D0;   // 266  0.774 
assign  ham[267] = 32'h624AE841;   // 267  0.768 
assign  ham[268] = 32'h617C53F9;   // 268  0.762 
assign  ham[269] = 32'h60ABF505;   // 269  0.755 
assign  ham[270] = 32'h5FD9D88E;   // 270  0.749 
assign  ham[271] = 32'h5F060BDA;   // 271  0.742 
assign  ham[272] = 32'h5E309C48;   // 272  0.736 
assign  ham[273] = 32'h5D599756;   // 273  0.729 
assign  ham[274] = 32'h5C810A96;   // 274  0.723 
assign  ham[275] = 32'h5BA703B8;   // 275  0.716 
assign  ham[276] = 32'h5ACB9080;   // 276  0.709 
assign  ham[277] = 32'h59EEBECC;   // 277  0.703 
assign  ham[278] = 32'h59109C8C;   // 278  0.696 
assign  ham[279] = 32'h583137CB;   // 279  0.689 
assign  ham[280] = 32'h57509EA3;   // 280  0.682 
assign  ham[281] = 32'h566EDF45;   // 281  0.675 
assign  ham[282] = 32'h558C07F3;   // 282  0.668 
assign  ham[283] = 32'h54A82701;   // 283  0.661 
assign  ham[284] = 32'h53C34AD4;   // 284  0.654 
assign  ham[285] = 32'h52DD81E1;   // 285  0.647 
assign  ham[286] = 32'h51F6DAAA;   // 286  0.640 
assign  ham[287] = 32'h510F63C2;   // 287  0.633 
assign  ham[288] = 32'h50272BC8;   // 288  0.626 
assign  ham[289] = 32'h4F3E4166;   // 289  0.619 
assign  ham[290] = 32'h4E54B354;   // 290  0.612 
assign  ham[291] = 32'h4D6A9050;   // 291  0.605 
assign  ham[292] = 32'h4C7FE726;   // 292  0.598 
assign  ham[293] = 32'h4B94C6A8;   // 293  0.590 
assign  ham[294] = 32'h4AA93DAF;   // 294  0.583 
assign  ham[295] = 32'h49BD5B1D;   // 295  0.576 
assign  ham[296] = 32'h48D12DD8;   // 296  0.569 
assign  ham[297] = 32'h47E4C4CB;   // 297  0.562 
assign  ham[298] = 32'h46F82EE4;   // 298  0.554 
assign  ham[299] = 32'h460B7B15;   // 299  0.547 
assign  ham[300] = 32'h451EB852;   // 300  0.540 
assign  ham[301] = 32'h4431F58F;   // 301  0.533 
assign  ham[302] = 32'h434541C0;   // 302  0.526 
assign  ham[303] = 32'h4258ABD9;   // 303  0.518 
assign  ham[304] = 32'h416C42CC;   // 304  0.511 
assign  ham[305] = 32'h40801586;   // 305  0.504 
assign  ham[306] = 32'h3F9432F4;   // 306  0.497 
assign  ham[307] = 32'h3EA8A9FC;   // 307  0.490 
assign  ham[308] = 32'h3DBD897E;   // 308  0.482 
assign  ham[309] = 32'h3CD2E054;   // 309  0.475 
assign  ham[310] = 32'h3BE8BD50;   // 310  0.468 
assign  ham[311] = 32'h3AFF2F3D;   // 311  0.461 
assign  ham[312] = 32'h3A1644DC;   // 312  0.454 
assign  ham[313] = 32'h392E0CE2;   // 313  0.447 
assign  ham[314] = 32'h384695FA;   // 314  0.440 
assign  ham[315] = 32'h375FEEC3;   // 315  0.433 
assign  ham[316] = 32'h367A25D0;   // 316  0.426 
assign  ham[317] = 32'h359549A2;   // 317  0.419 
assign  ham[318] = 32'h34B168B0;   // 318  0.412 
assign  ham[319] = 32'h33CE915E;   // 319  0.405 
assign  ham[320] = 32'h32ECD200;   // 320  0.398 
assign  ham[321] = 32'h320C38D9;   // 321  0.391 
assign  ham[322] = 32'h312CD417;   // 322  0.384 
assign  ham[323] = 32'h304EB1D8;   // 323  0.377 
assign  ham[324] = 32'h2F71E024;   // 324  0.371 
assign  ham[325] = 32'h2E966CEC;   // 325  0.364 
assign  ham[326] = 32'h2DBC660D;   // 326  0.357 
assign  ham[327] = 32'h2CE3D94E;   // 327  0.351 
assign  ham[328] = 32'h2C0CD45B;   // 328  0.344 
assign  ham[329] = 32'h2B3764CA;   // 329  0.338 
assign  ham[330] = 32'h2A639816;   // 330  0.331 
assign  ham[331] = 32'h29917B9F;   // 331  0.325 
assign  ham[332] = 32'h28C11CAB;   // 332  0.318 
assign  ham[333] = 32'h27F28863;   // 333  0.312 
assign  ham[334] = 32'h2725CBD4;   // 334  0.306 
assign  ham[335] = 32'h265AF3ED;   // 335  0.300 
assign  ham[336] = 32'h25920D7D;   // 336  0.294 
assign  ham[337] = 32'h24CB2535;   // 337  0.287 
assign  ham[338] = 32'h240647A5;   // 338  0.281 
assign  ham[339] = 32'h2343813D;   // 339  0.275 
assign  ham[340] = 32'h2282DE4A;   // 340  0.270 
assign  ham[341] = 32'h21C46AF7;   // 341  0.264 
assign  ham[342] = 32'h2108334B;   // 342  0.258 
assign  ham[343] = 32'h204E432B;   // 343  0.252 
assign  ham[344] = 32'h1F96A654;   // 344  0.247 
assign  ham[345] = 32'h1EE16860;   // 345  0.241 
assign  ham[346] = 32'h1E2E94C2;   // 346  0.236 
assign  ham[347] = 32'h1D7E36C5;   // 347  0.230 
assign  ham[348] = 32'h1CD0598C;   // 348  0.225 
assign  ham[349] = 32'h1C250814;   // 349  0.220 
assign  ham[350] = 32'h1B7C4D2F;   // 350  0.215 
assign  ham[351] = 32'h1AD63384;   // 351  0.210 
assign  ham[352] = 32'h1A32C593;   // 352  0.205 
assign  ham[353] = 32'h19920DAC;   // 353  0.200 
assign  ham[354] = 32'h18F415F8;   // 354  0.195 
assign  ham[355] = 32'h1858E871;   // 355  0.190 
assign  ham[356] = 32'h17C08EE3;   // 356  0.186 
assign  ham[357] = 32'h172B12EE;   // 357  0.181 
assign  ham[358] = 32'h16987E04;   // 358  0.177 
assign  ham[359] = 32'h1608D967;   // 359  0.172 
assign  ham[360] = 32'h157C2E29;   // 360  0.168 
assign  ham[361] = 32'h14F2852E;   // 361  0.164 
assign  ham[362] = 32'h146BE726;   // 362  0.160 
assign  ham[363] = 32'h13E85C93;   // 363  0.156 
assign  ham[364] = 32'h1367EDC4;   // 364  0.152 
assign  ham[365] = 32'h12EAA2D5;   // 365  0.148 
assign  ham[366] = 32'h127083B1;   // 366  0.144 
assign  ham[367] = 32'h11F9980E;   // 367  0.140 
assign  ham[368] = 32'h1185E770;   // 368  0.137 
assign  ham[369] = 32'h11157924;   // 369  0.133 
assign  ham[370] = 32'h10A85445;   // 370  0.130 
assign  ham[371] = 32'h103E7FB8;   // 371  0.127 
assign  ham[372] = 32'h0FD8022C;   // 372  0.124 
assign  ham[373] = 32'h0F74E21B;   // 373  0.121 
assign  ham[374] = 32'h0F1525C6;   // 374  0.118 
assign  ham[375] = 32'h0EB8D33B;   // 375  0.115 
assign  ham[376] = 32'h0E5FF04E;   // 376  0.112 
assign  ham[377] = 32'h0E0A829C;   // 377  0.110 
assign  ham[378] = 32'h0DB88F8C;   // 378  0.107 
assign  ham[379] = 32'h0D6A1C49;   // 379  0.105 
assign  ham[380] = 32'h0D1F2DC8;   // 380  0.103 
assign  ham[381] = 32'h0CD7C8C6;   // 381  0.100 
assign  ham[382] = 32'h0C93F1C4;   // 382  0.098 
assign  ham[383] = 32'h0C53AD0B;   // 383  0.096 
assign  ham[384] = 32'h0C16FEAC;   // 384  0.094 
assign  ham[385] = 32'h0BDDEA7A;   // 385  0.093 
assign  ham[386] = 32'h0BA87411;   // 386  0.091 
assign  ham[387] = 32'h0B769ED2;   // 387  0.090 
assign  ham[388] = 32'h0B486DE2;   // 388  0.088 
assign  ham[389] = 32'h0B1DE42C;   // 389  0.087 
assign  ham[390] = 32'h0AF70460;   // 390  0.086 
assign  ham[391] = 32'h0AD3D0F3;   // 391  0.085 
assign  ham[392] = 32'h0AB44C1D;   // 392  0.084 
assign  ham[393] = 32'h0A9877DD;   // 393  0.083 
assign  ham[394] = 32'h0A8055F4;   // 394  0.082 
assign  ham[395] = 32'h0A6BE7E9;   // 395  0.081 
assign  ham[396] = 32'h0A5B2F05;   // 396  0.081 
assign  ham[397] = 32'h0A4E2C59;   // 397  0.081 
assign  ham[398] = 32'h0A44E0B4;   // 398  0.080 
assign  ham[399] = 32'h0A3F4CB0;   // 399  0.080 

endmodule